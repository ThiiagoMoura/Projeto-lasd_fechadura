module Memoria_Instrucao (A, RD);

input [7:0] A;

output reg [31:0] RD;


always @(*)begin
	case(A)
		8'b00000000: RD = 32'b_001000_00000_00001_00000_00000_000011; 
		8'b00000001: RD = 32'b_001000_00000_00010_00000_00000_001001;
		8'b00000010: RD = 32'b_000000_00001_00010_00010_00000_100000;
		8'b00000011: RD = 32'b_000000_00001_00010_00011_00000_100100;
		8'b00000100: RD = 32'b_000000_00001_00010_00100_00000_100101;
		8'b00000101: RD = 32'b001000_00001_00000_00000_00000_000010;
		default:     RD = 32'b001000_00000_00000_00000_00000_000000;
					
	endcase
end



endmodule
